module top (output rgb0_g);
   (* KEEP, DONT_TOUCH *)
   LUT2 #( .INIT(4'b0) ) lut ( .O(rgb0_g));

endmodule
