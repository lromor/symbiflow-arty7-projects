module top (output rgb0_g);
   reg t = 1'b0;
endmodule
